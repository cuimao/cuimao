#include "uvm.sv"
